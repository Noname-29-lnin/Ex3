task automatic Simulus_data();
    begin
        
    end
endtask //automatic