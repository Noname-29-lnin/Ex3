task Display_Data();
    begin
        $display("Output data \n");
    end
endtask
