class transaction_driver;

endclass
